module shifter(
		input  [31:0] A,
		input  [ 7:0] BY,	// How many bits it needs to shifted by 
		
		output [31:0] OUT
	);
	
endmodule 